module proc(i_clk, i_rst);
    input    i_clk, i_rst;

    wire [31:0] pc, pc_inc, pc_next, pc_jump, val_reg0, val_reg1,
                         ram_addr, ram_out, wb_val_alu, wb_val, alu_out;
    wire [15:0] ir;
    wire [ 4:0] reg0, reg1, wb_reg;
    wire [ 3:0] inst, alu_action;
    wire [ 1:0] fmt, ram_action;
    wire        do_jump;
 
    pc        pc_(.i_clk(i_clk),
                  .i_rst(i_rst),
                  .i_pc(pc_next),
                  .o_pc(pc),
                  .o_pc_inc(pc_inc));
 
    /* TODO: there should be no ROM, instead only one RAM module */
    rom        rom(.i_addr(pc),
                   .o_data(ir));

    dispatcher dispatcher(.i_ir(ir),
                          .o_fmt(fmt),
                          .o_inst(inst),
                          .o_reg0(reg0),
                          .o_reg1(reg1));

    regf        regf(.i_clk(i_clk),
                     .i_reg0(reg0),
                     .i_reg1(reg1),
                     .i_wb_reg(wb_reg),
                     .i_wb_val(wb_val),
                     .o_reg0(val_reg0),
                     .o_reg1(val_reg1));

    control     control(.i_clk(i_clk),
                        .i_inst(inst),
                        .i_reg0(reg0),
                        .i_reg1(reg1),
                        .i_val_reg0(val_reg0),
                        .i_val_reg1(val_reg1),
                        .i_pc_inc(pc_inc),
                        .i_alu_out(alu_out),
                        .o_ram_action(ram_action),
                        .o_ram_addr(ram_addr),
                        .o_do_jump(do_jump),
                        .o_alu_action(alu_action),
                        .o_wb_reg(wb_reg),
                        .o_wb_val(wb_val));

    alu_total   alu(.i_reg0(val_reg0),
                    .i_reg1(val_reg1),
                    .i_alu_action(alu_action),
                    .i_fmt(fmt),
                    .o_alu_out(alu_out));

    ram      ram(.i_clk(i_clk),
                 .i_action(ram_action),
                 .i_addr(ram_addr),
                 .i_val(val_reg0),
                 .o_val(ram_out));

   assign pc_jump = val_reg1;
   assign pc_next = (do_jump ? pc_inc : pc_jump);

endmodule

